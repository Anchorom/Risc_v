module ctrl (


);









endmodule
